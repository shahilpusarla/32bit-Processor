// Datamemory module
module memory_16_32d(data,data2,addr,ins1,clk);
output [31:0] data;
input  [31:0] addr,data2;
input [5:0]ins1;
input clk;
reg [31:0] data;
reg [31:0] memdata [255:0];

initial 
	begin
	memdata[0] = 32'b00000000000000000000000000000000;
	memdata[1] = 32'b00000000000000000000000000000001;
	memdata[2] = 32'b00000000000000000000000000000010;
	memdata[3] = 32'b00000000000000000000000000000011;
	memdata[4] = 32'b00000000000000000000000000000100;
	memdata[5] = 32'b00000000000000000000000000000101;
	memdata[6] = 32'b00000000000000000000000000000110;
	memdata[7] = 32'b00000000000000000000000000000111;
	memdata[8] = 32'b00000000000000000000000000001000;
	memdata[9] = 32'b00000000000000000000000000001001;
	memdata[10] = 32'b00000000000000000000000000001010;
	memdata[11] = 32'b00000000000000000000000000001011;
	memdata[12] = 32'b00000000000000000000000000001100;
	memdata[13] = 32'b00000000000000000000000000001101;
	memdata[14] = 32'b00000000000000000000000000001110;
	memdata[15] = 32'b00000000000000000000000000001111;
	memdata[16] = 32'b00000000000000000000000000010000;
	memdata[17] = 32'b00000000000000000000000000010001;
	memdata[18] = 32'b00000000000000000000000000100000;
	memdata[19] = 32'b00000000000000000000000000100000;
	memdata[20] = 32'b00000000000000000000000001000000;
	memdata[21] = 32'b00000000000000000000000001000000;
	memdata[22] = 32'b00000000000000000000000010000000;
	memdata[23] = 32'b00000000000000000000000010000000;
	memdata[24] = 32'b00000000000000000000000100000000;
	memdata[25] = 32'b00000000000000000000000100000000;
	memdata[26] = 32'b00000000000000000000000100000000;
	memdata[27] = 32'b00000000000000000000000100000000;
	memdata[28] = 32'b00000000000000000000011000000000;
	memdata[29] = 32'b00000000000000000000110000000000;
	memdata[30] = 32'b00000000000000000000000000000000;
	memdata[31] = 32'b00000000000000000000001000000000;
	memdata[32] = 32'b00000000000000000000110000000000;	
	memdata[33] = 32'b00000000000000000000001010000000;
	memdata[34] = 32'b00000000000000000000011100000000;
	memdata[35] = 32'b00000000000000000000001111000000;
	memdata[36] = 32'b00000000000000000000111110000000;
	memdata[37] = 32'b00000000000000000000000010000000;
	memdata[38] = 32'b00000000000000000010000000000000;
	memdata[39] = 32'b00000000000000000010100000000000;
	memdata[40] = 32'b00000000000000000000100000000000;
	memdata[41] = 32'b00000000000000000000010000000000;
	memdata[42] = 32'b00000000000000000000100000000000;
	memdata[43] = 32'b00000000000000000001000000000000;
	memdata[44] = 32'b00000000000000000000010000000000;
	memdata[45] = 32'b00000000000000000000010000000000;
	memdata[46] = 32'b00000000000000000000100000000000;
	memdata[47] = 32'b00000000000000000000100000000000;
	memdata[48] = 32'b00000000000000000000110000000000;
	memdata[49] = 32'b00000000000000000000010000000000;
	memdata[50] = 32'b00000000000000000000011000000000;
	memdata[51] = 32'b00000000000000000000011000000000;
	memdata[52] = 32'b00000000000000000000001000000000;
	memdata[53] = 32'b00000000000000000000000100000000;
	memdata[54] = 32'b00000000000000000000000000000000;
	memdata[55] = 32'b00000000000000000000000100000000;
	memdata[56] = 32'b00000000000000000000000100000000;
	memdata[57] = 32'b00000000000000000000001000000000;
	memdata[58] = 32'b00000000000000000000100000000000;
	memdata[59] = 32'b00000000000000000000100000000000;
	memdata[60] = 32'b00000000000000000001000000000000;
	memdata[61] = 32'b00000000000000000010000000000000;
	memdata[62] = 32'b00000000000000000010000000000000;
	memdata[63] = 32'b00000000000000000010000000000000;
	memdata[64] = 32'b00000000000000000010000000000000;
	memdata[65] = 32'b00000000000000001000000000000000;
	memdata[66] = 32'b00000000000000010000000000000000;
	memdata[67] = 32'b00000000000000100000000000000000;
	memdata[68] = 32'b00000000000000100000000000000000;
	memdata[69] = 32'b00000000000000100000000000000000;
	memdata[70] = 32'b00000000000000110000000000000000;
	memdata[71] = 32'b00000000000000010000000000000000;
	memdata[72] = 32'b00000000000000010000000000000000;
	memdata[73] = 32'b00000000000000000000000000000000;
	memdata[74] = 32'b00000000000000000000000000000000;
	memdata[75] = 32'b00000000000000000000000000000000;
	memdata[76] = 32'b00000000000000000000000000000000;
	memdata[77] = 32'b00000000000000000000000000000000;
	memdata[78] = 32'b00000000000000000000000000000000;
	memdata[79] = 32'b00000000000000000000000000000000;
	memdata[80] = 32'b00000000000000000000000000000000;
	memdata[81] = 32'b00000000000000000000000000000000;
	memdata[82] = 32'b00000000000000000000000000000000;
	memdata[83] = 32'b00000000000000000000000000000000;
	memdata[84] = 32'b00000000000000000000000000000000;
	memdata[85] = 32'b00000000000000000000000000000000;
	memdata[86] = 32'b00000000000000000000000000000000;
	memdata[87] = 32'b00000000000000000000000000000000;
	memdata[88] = 32'b00000000000000000000000000000000;
	memdata[89] = 32'b00000000000000000000000000000000;
	memdata[90] = 32'b00000000000000000000000000000000;
	memdata[91] = 32'b00000000000000000000000000000000;
	memdata[92] = 32'b00000000000000000000000000000000;
	memdata[93] = 32'b00000000000000000000000000000000;
	memdata[94] = 32'b00000000000000000000000000000000;
	memdata[95] = 32'b00000000000000000000000000000000;
	memdata[96] = 32'b00000000000000000000000000000000;
	memdata[97] = 32'b00000000000000000000000000000000;	
	memdata[98] = 32'b00000000000000000000000000000000;
	memdata[99] = 32'b00000000000000000000000000000000;
	memdata[100] = 32'b00000000000000000000000000000000;
	memdata[101] = 32'b00000000000000000000000000000000;
	memdata[102] = 32'b00000000000000000000000000000000;
	memdata[103] = 32'b00000000000000000000000000000000;
	memdata[104] = 32'b00000000000000000000000000000000;
	memdata[105] = 32'b00000000000000000000000000000000;
	memdata[106] = 32'b00000000000000000000000000000000;
	memdata[107] = 32'b00000000000000000000000000000000;
	memdata[108] = 32'b00000000000000000000000000000000;
	memdata[109] = 32'b00000000000000000000000000000000;
	memdata[110] = 32'b00000000000000000000000000000000;
	memdata[111] = 32'b00000000000000000000000000000000;
	memdata[112] = 32'b00000000000000000000000000000000;
	memdata[113] = 32'b00000000000000000000000000000000;
	memdata[114] = 32'b00000000000000000000000000000000;
	memdata[115] = 32'b00000000000000000000000000000000;
	memdata[116] = 32'b00000000000000000000000000000000;
	memdata[117] = 32'b00000000000000000000000000000000;
	memdata[118] = 32'b00000000000000000000000000000000;
	memdata[119] = 32'b00000000000000000000000000000000;
	memdata[120] = 32'b00000000000000000000000000000000;
	memdata[121] = 32'b00000000000000000000000000000000;
	memdata[122] = 32'b00000000000000000000000000000000;
	memdata[123] = 32'b00000000000000000000000000000000;
	memdata[124] = 32'b00000000000000000000000000000000;
	memdata[125] = 32'b00000000000000000000000000000000;
	memdata[126] = 32'b00000000000000000000000000000000;
	memdata[127] = 32'b00000000000000000000000000000000;
	memdata[128] = 32'b00000000000000000000000000000000;
	memdata[129] = 32'b00000000000000000000000000000000;	
	end

always @(clk)
	begin
	if(ins1==6'b100011)
		data = memdata[addr];
	else if(ins1 == 6'b000001)
		data = addr; 
	if(ins1==6'b101011)
		memdata[addr] = data2;
	end
endmodule


//Instruction Memory Module

module memory_16_32i(data1,data2,data3,data4,ins4_rd,ins4alu,da,addr,clk);
output [5:0] data1;
output [4:0] data2,data3;
output [15:0] data4;
output [5:0]ins4alu;
output [4:0]ins4_rd;
output [31:0]da;
input  [15:0] addr;
input clk;
reg [5:0] data1,ins4alu;
reg [15:0] data4;
reg [31:0]da;
reg [4:0] data3,data2,ins4_rd;
reg [5:0] memdata1 [127:0];
reg [15:0] memdata4 [127:0];
reg [4:0] memdata2 [127:0];
reg [4:0] memdata3 [127:0];
initial 
	begin
	memdata1[0] = 6'b100011;
	memdata2[0] = 5'b00000;
	memdata3[0] = 5'b00001;
	memdata4[0] =16'b0000000000100000;
	memdata1[1] = 6'b100011;
	memdata2[1] = 5'b00001;
	memdata3[1] = 5'b00011;
	memdata4[1] =16'b0000000000100100;
        memdata1[2] = 6'b100011;
	memdata2[2] = 5'b00101;
	memdata3[2] = 5'b00011;
	memdata4[2] =16'b0000000001100000;
	memdata1[3] = 6'b000001;
	memdata2[3] = 5'b00001;
	memdata3[3] = 5'b00111;
	memdata4[3] =16'b0000000000100000;
	memdata1[4] = 6'b000001;
	memdata2[4] = 5'b00010;
	memdata3[4] = 5'b00111;
	memdata4[4] =16'b0000000000100000;
	memdata1[5] = 6'b000001;
	memdata2[5] = 5'b00011;
	memdata3[5] = 5'b00001;
	memdata4[5] =16'b0000000000100010;
	memdata1[6] = 6'b000001;
	memdata2[6] = 5'b00001;
	memdata3[6] = 5'b00011;
	memdata4[6] =16'b0000000000100010;
	memdata1[7] = 6'b000001;
	memdata2[7] = 5'b00001;
	memdata3[7] = 5'b00010;
	memdata4[7] =16'b0000000000100100;
	memdata1[8] = 6'b000001;
	memdata2[8] = 5'b00010;
	memdata3[8] = 5'b00011;
	memdata4[8] =16'b0000000000100100;
	memdata1[9] = 6'b000001;
	memdata2[9] = 5'b00001;
	memdata3[9] = 5'b00010;
	memdata4[9] =16'b0000000000100101;
	memdata1[10] = 6'b000001;
	memdata2[10] = 5'b00010;
	memdata3[10] = 5'b00010;
	memdata4[10] =16'b000000000100101;
	memdata1[11] = 6'b101011;
	memdata2[11] = 5'b00000;
	memdata3[11] = 5'b00000;
	memdata4[11] =16'b0000000000101011;
	memdata1[12] = 6'b101011;
	memdata2[12] = 5'b00001;
	memdata3[12] = 5'b00000;
	memdata4[12] =16'b0000000000101011;
	memdata1[13] = 6'b000010;
	memdata2[13] = 5'b00001;
	memdata3[13] = 5'b00001;
	memdata4[13] =16'b0000000000000011;
	memdata1[14] = 6'b000001;
	memdata2[14] = 5'b00001;
	memdata3[14] = 5'b00000;
	memdata4[14] =16'b0000000000100000;
	memdata1[15] = 6'b000001;
	memdata2[15] = 5'b00001;
	memdata3[15] = 5'b00000;
	memdata4[15] =16'b0000000000100000;
	memdata1[16] = 6'b000001;
	memdata2[16] = 5'b00001;
	memdata3[16] = 5'b00011;
	memdata4[16] =16'b0000000000100000;
	memdata1[17] = 6'b000001;
	memdata2[17] = 5'b00001;
	memdata3[17] = 5'b00011;
	memdata4[17] =16'b0000000000100000;
	memdata1[18] = 6'b000001;
	memdata2[18] = 5'b00001;
	memdata3[18] = 5'b00011;
	memdata4[18] =16'b0000000000100000;
	end

always @(posedge clk)
	begin
		data1 = memdata1[addr];
		data2 = memdata2[addr];
		data3 = memdata3[addr];
		data4 = memdata4[addr];
		ins4_rd[4] = data4[15];
		ins4_rd[3] = data4[14];
		ins4_rd[2] = data4[13];
		ins4_rd[1] = data4[12];
		ins4_rd[0] = data4[11];
		ins4alu[0] = data4[0];
		ins4alu[1] = data4[1];
		ins4alu[2] = data4[2];
		ins4alu[3] = data4[3];
		ins4alu[4] = data4[4];
		ins4alu[5] = data4[5];
		da = data4;
	end
endmodule


//clk Module

module clock(out);
output out;
reg out;

initial begin
	out = 1'b0;
end

always 
	begin
		out = #1 ~out;
	end
endmodule

//Counter Module
module counter(out,en,reset,ins4,ins1,clk);
output [15:0] out;
reg    [15:0] out;
input [15:0]ins4;
input [5:0]ins1;
input  en,reset,clk;
always @(posedge clk or reset)
begin
	if(reset == 1'b1)
	begin
		out = 16'b0000000000000000;
	end
	else if(en == 1'b1 && ins1 != 6'b000010)
	begin
		out = out + 1;
	end
	else if(en == 1'b1 && ins1 == 6'b000010)
		begin
		out = out + ins4;
		end 
end
endmodule

//Register File Module

module memory_16_32r(data1,data2,ins2,ins3,ins4_rd,ins1,medi,clk);
output [31:0] data1,data2;
input  [4:0] ins2,ins3;
input [4:0]ins4_rd;
input [5:0]ins1;
input clk;
input [31:0]medi;
reg [31:0] data1,data2;
reg [31:0] memdata [31:0];
initial begin
	memdata[0] = 32'b00000000000000000000000000000001;
	memdata[1] = 32'b00000000000000000000000000000001;
	memdata[2] = 32'b00000000000000000000000000000010;
	memdata[3] = 32'b00000000000000000000000000000011;
	memdata[4] = 32'b00000000000000000000000000000011;
	memdata[5] = 32'b00000000000000000000000000000010;
	memdata[6] = 32'b00000000000000000000000000000001;
	memdata[7] = 32'b00000000000000000000000000000011;
	memdata[8] = 32'b00000000000000000000000000000010;
	memdata[9] = 32'b00000000000000000000000000000001;
	memdata[10] = 32'b00000000000000000000000000000011;
	memdata[11] = 32'b00000000000000000000000000000111;
	memdata[12] = 32'b00000000000000000000000000001011;
	memdata[13] = 32'b00000000000000000000000000001001;
	memdata[14] = 32'b00000000000000000000000000001101;
	memdata[15] = 32'b00000000000000000000000000000001;
	memdata[16] = 32'b00000000000000000000000000000001;
	memdata[17] = 32'b00000000000000000000000000000001;
	memdata[18] = 32'b00000000000000000000000000000001;
	memdata[19] = 32'b00000000000000000000000000000001;
	memdata[20] = 32'b00000000000000000000000000000000;
	memdata[21] = 32'b00000000000000000000000000000000;
	memdata[22] = 32'b00000000000000000000000000000000;
	memdata[23] = 32'b00000000000000000000000000000000;
	memdata[24] = 32'b00000000000000000000000000000000;
	memdata[25] = 32'b00000000000000000000000000000000;
	memdata[26] = 32'b00000000000000000000000000000000;
	memdata[27] = 32'b00000000000000000000000000000000;
	memdata[28] = 32'b00000000000000000000000000000000;
	memdata[29] = 32'b00000000000000000000000000000000;
	memdata[30] = 32'b00000000000000000000000000000000;
	memdata[31] = 32'b00000000000000000000000000000000;
end
always @(posedge clk)
	begin
		data1 = memdata[ins2];
		data2 = memdata[ins3];
	end
always @(posedge clk)
begin
if(ins1==6'b000001 || ins1==6'b100011)
memdata[ins4_rd] = medi;
end
endmodule


//ALU module

module Alu(data,data1,data2,data3,ins4,ins1,clk);
input [5:0]ins4;
input [5:0]ins1;
output [31:0]data;
reg [31:0]data;
input [31:0]data1,data2,data3;
input clk;
always @(negedge clk)
begin
if(ins1==6'b100011 || ins1==6'b101011)
begin
data=data1+data2;
end
else if(ins1==6'b000001 && ins4[0]==0 && ins4[1]==0 && ins4[2]==0 && ins4[3]==0 && ins4[4]==0 && ins4[5]==1)
begin
data=data1 + data3;
end
else if(ins1==6'b000001 && ins4[0]==0 && ins4[1]==0 && ins4[2]==1 && ins4[3]==0 && ins4[4]==0 && ins4[5]==1)
begin
data=data1 & data3;
end
else if(ins1==6'b000001 && ins4[0]==1 && ins4[1]==0 && ins4[2]==1 && ins4[3]==0 && ins4[4]==0 && ins4[5]==1)
begin
data=data1 | data3;
end
else if(ins1==6'b000001 && ins4[0]==0 && ins4[1]==1 && ins4[2]==0 && ins4[3]==0 && ins4[4]==0 && ins4[5]==1)
begin
data=data1-data3;
end
else if(ins1 == 6'b000010)
begin
data=data1-data3;
end
end
endmodule

//Test Bench

module TB;
reg en,reset;
wire [5:0]ins1;
wire [4:0]ins2,ins3;
wire [15:0]ins4;
wire [4:0]ins4_rd;
wire [5:0]ins4alu;
wire [15:0]addr;
wire [31:0]da,data1,data2,data,datamemory;
reg [31:0]mediator;
clock clk01(clk);
counter c(addr,en,reset,ins4,ins1,clk);

memory_16_32i m1(ins1,ins2,ins3,ins4,ins4_rd,ins4alu,da,addr,clk);
memory_16_32r m3(data1,data2,ins2,ins3,ins4_rd,ins1,mediator,clk);
Alu A1(data,data1,da,data2,ins4alu,ins1,clk);
memory_16_32d m4(datamemory,data2,data,ins1,clk);

initial begin
$monitor("destination reg value,rt in load case and rd in other operations case except beq and store =%b \n Address to access in datamemory for load/store and operation value in other operations=%b \nopcode=%brs=%brt=%baddr=%b rs-data=%b rt-data=%b clk=%b pc=%d", datamemory,data,ins1,ins2,ins3,ins4,data1,data2,clk,addr);
reset=1'b1;
#1 en=1'b1;
reset = 1'b0;
#30
$finish;
end
always @(data)
begin
if(ins1==6'b000001)
mediator=datamemory;
else if(ins1==6'b100011)
mediator=datamemory;
end 
endmodule
